module lab1_AND_GATE
(
input  A,
input B,
output Y
);
assign Y=A&B;
endmodule
